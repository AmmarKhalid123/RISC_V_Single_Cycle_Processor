module Instruction_Memory
(
  input [63:0]Instr_Addr,
  output reg [31:0]Instruction
);

reg [7:0]regs[95:0];

initial
begin



        regs[0] = 8'b00010011; 
        regs[1] = 8'b00001011; 
        regs[2] = 8'b00000000; 
        regs[3] = 8'b00000000; 

        regs[4] = 8'b00010011; 
        regs[5] = 8'b00000101; 
        regs[6] = 8'b01010000; 
        regs[7] = 8'b00000000; 

        regs[8] = 8'b00010011; 
        regs[9] = 8'b00000001; 
        regs[10] = 8'b00000000; 
        regs[11] = 8'b00000000; 

        regs[12] = 8'b10010011; 
        regs[13] = 8'b00000001; 
        regs[14] = 8'b00000000; 
        regs[15] = 8'b00000000; 
          
        regs[16] = 8'b10110011; 
        regs[17] = 8'b00001011; 
        regs[18] = 8'b01100000; 
        regs[19] = 8'b00000001; 

        regs[20] = 8'b01100011; 
        regs[21] = 8'b00000110; 
        regs[22] = 8'b10101011; 
        regs[23] = 8'b00000100; 

        regs[24] = 8'b00000011; 
        regs[25] = 8'b00110011; 
        regs[26] = 8'b00000001; 
        regs[27] = 8'b00000000; 

        regs[28] = 8'b00000011; 
        regs[29] = 8'b10110010; 
        regs[30] = 8'b00000001; 
        regs[31] = 8'b00000000;

        regs[32] = 8'b01100011; 
        regs[33] = 8'b01001110; 
        regs[34] = 8'b01000011; 
        regs[35] = 8'b00000000; 

        regs[36] = 8'b10010011; 
        regs[37] = 8'b10001011; 
        regs[38] = 8'b00011011; 
        regs[39] = 8'b00000000; 

        regs[40] = 8'b00010011; 
        regs[41] = 8'b00010001; 
        regs[42] = 8'b00111011; 
        regs[43] = 8'b00000000; 

        regs[44] = 8'b10010011; 
        regs[45] = 8'b10010001; 
        regs[46] = 8'b00111011; 
        regs[47] = 8'b00000000; 

        regs[48] = 8'b11100011; 
        regs[49] = 8'b10010100; 
        regs[50] = 8'b10101011; 
        regs[51] = 8'b11111110; 

        regs[52] = 8'b00010011; 
        regs[53] = 8'b00001011; 
        regs[54] = 8'b00011011; 
        regs[55] = 8'b00000000; 

        regs[56] = 8'b11100011; 
        regs[57] = 8'b10001100; 
        regs[58] = 8'b10101011; 
        regs[59] = 8'b11111100; 

        regs[60] = 8'b10110011; 
        regs[61] = 8'b00000010; 
        regs[62] = 8'b01100000; 
        regs[63] = 8'b00000000; 

        regs[64] = 8'b00100011; 
        regs[65] = 8'b00110000; 
        regs[66] = 8'b01000001; 
        regs[67] = 8'b00000000; 

        regs[68] = 8'b00100011; 
        regs[69] = 8'b10110000; 
        regs[70] = 8'b01010001; 
        regs[71] = 8'b00000000; 

        regs[72] = 8'b10010011; 
        regs[73] = 8'b10001011; 
        regs[74] = 8'b00011011; 
        regs[75] = 8'b00000000;

        regs[76] = 8'b00010011; 
        regs[77] = 8'b00010001; 
        regs[78] = 8'b00111011; 
        regs[79] = 8'b00000000;

        regs[80] = 8'b10010011; 
        regs[81] = 8'b10010001; 
        regs[82] = 8'b00111011; 
        regs[83] = 8'b00000000;

        regs[84] = 8'b11100011; 
        regs[85] = 8'b10010010; 
        regs[86] = 8'b10101011; 
        regs[87] = 8'b11111100;

        regs[88] = 8'b00010011; 
        regs[89] = 8'b00001011; 
        regs[90] = 8'b00011011; 
        regs[91] = 8'b00000000;

        regs[92] = 8'b11100011; 
        regs[93] = 8'b10001010; 
        regs[94] = 8'b10101011; 
        regs[95] = 8'b11111010;

end

always @ (Instr_Addr)
begin
  Instruction = {regs[Instr_Addr + 2'b11], regs[Instr_Addr + 2'b10], regs[Instr_Addr + 1'b1], regs[Instr_Addr]};
end

endmodule