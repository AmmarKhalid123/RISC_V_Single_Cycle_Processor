module ALU_Control
(
  input [1:0]ALUOp,
  input [3:0]Funct,
  output reg [3:0]Operation
);

always @ (ALUOp, Funct)
begin
  if (ALUOp == 2'b00)
    begin
      case(Funct)
        4'b0001 : Operation = 4'b0100; //slli
        default : Operation = 4'b0010;
      endcase
    end
  if (ALUOp == 2'b01)
    begin
      case({Funct})
        4'b0000 : Operation = 4'b0110; //beq
	4'b0001 : Operation = 4'b0011; //bne
	4'b0100 : Operation = 4'b0111; //blt
      endcase
    end
  if (ALUOp == 2'b10)
    begin
      if (Funct == 4'b0000)
	begin
          Operation = 4'b0010;
	end
      if (Funct == 4'b1000)
	begin
          Operation <= 4'b0110;
	end
      if (Funct == 4'b0111)
	begin
          Operation = 4'b0000;
	end
      if (Funct == 4'b0110)
        begin
	  Operation = 4'b0001;
	end
    end
end

endmodule